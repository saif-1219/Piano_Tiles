`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 05/10/2023 02:58:25 PM
// Design Name: 
// Module Name: top_of_the_tops
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


//module top_of_the_tops(
//input clk,
//input button_1,
//input button_2,
//input button_3,
//input button_4,
//input start_button,
//input x,
//input y,
//input [3:0] state,
//input st_change,
//input video_on,
//output [3:0] red,
//output [3:0] green,
//output [3:0] blue
//    );
//reg [1:0] game_state = 0;

//if (game_state==0) begin
//    pix_gen_menu menu(clk,x,y,start_button,video_on,red,green,blue,game_state);
//    end

 
//endmodule
